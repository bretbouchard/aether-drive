* SPICE Netlist for Test LED Circuit
* Created: 2026-01-16
* Purpose: [Describe circuit purpose]

* ============================================================
* POWER SUPPLY
* ============================================================
VCC 1 0 DC 5.0

* ============================================================
* CIRCUIT DESCRIPTION
* ============================================================
[Add your circuit here]

* ============================================================
* SIMULATION
* ============================================================
.TRAN 10u 10m
.PRINT V(1) V(2)
.END
